library ieee;
use ieee.std_logic_1164.all;


entity BW_XOR is
  generic(
    n: integer := 6
  );
	port(
		grygorczuk_xor_1, grygorczuk_xor_2: in std_logic_vector(n-1 DOWNTO 0);
		grygorczuk_output_xor: out std_logic_vector(n-1 DOWNTO 0)
	);
end BW_XOR;

architecture BW_XOR_LOGIC of BW_XOR is

begin

XOR_LOOP: for i in 0 to n-1 generate
  grygorczuk_output_xor(i) <= grygorczuk_xor_1(i) xor grygorczuk_xor_2(i);
end generate;
  
end BW_XOR_LOGIC;